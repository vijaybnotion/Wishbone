-- See the file "LICENSE" for the full license governing this code. --

package lt16soc_utils is

	--insert utility component and function declarations

end lt16soc_utils;

package body lt16soc_utils is

	--insert utility function bodies

end lt16soc_utils;

